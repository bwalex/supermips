`define clogb2(n) $clog2(n)